module Video (
    input i_clk,
    input logic [9:0] i_pixel_x,
    input logic [8:0] i_pixel_y,
    input logic [1:0] i_state,
    output logic [15:0] o_color
);

    // wire setup
    logic [12:0] w_tile_addr;
    assign w_tile_addr = {i_pixel_y[8:3], i_pixel_x[9:3]};

    logic [2:0] w_tile_x, w_tile_y;
    assign w_tile_x = i_pixel_x[2:0];
    assign w_tile_y = i_pixel_y[2:0];

    // palette init
    logic [15:0] color [0:1];
    assign color[0] = (i_pixel_x[3] ^ i_pixel_y[3]) ? 16'hF100 : 16'h0000;
    assign color[1] = 16'hFFFF;

    // Tile index memory
    logic [7:0] w_tile_index;
    memory8k tilemap_inst (
        .i_clk(i_clk),
        .wen(1'b0),
        .ren(1'b1),
        .waddr(13'b0),
        .raddr(w_tile_addr),
        .wdata(8'b0),
        .rdata(w_tile_index)
    );

    logic [10:0] w_rom_addr;
    assign w_rom_addr = {w_tile_index, i_pixel_y[2:0]};
    logic [7:0] current_line;
    memory2k tilerom_inst (
        .i_clk(i_clk),
        .wen(1'b0),
        .ren(1'b1),
        .waddr(11'b0),
        .raddr(w_rom_addr),
        .wdata(8'b0),
        .rdata(current_line)
    );

    always_ff @(posedge i_clk) begin
       o_color <= color[current_line[~i_pixel_x[2:0]]];
    end
    
endmodule